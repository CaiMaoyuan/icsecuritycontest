package ariane_soc_pkg;        

        //HMAC key 
        localparam logic [31:0] HMACKey_3    =  17;
        localparam HMACKey_2    =  18;
        localparam HMACKey_1    =  19;
        localparam HMACKey_0    =  20;
endpackage
